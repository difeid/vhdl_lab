33&Файл зашифрован с помощью CryptCode.py 
33&Хфнкцжисѕє'&Иё&цжчюоъцфижсо&рфк2&фчшжсфчђ&хфтлуѕшђ&тлчшжто&хжцщ&зщри

ryhxgx&OKKKA
{ok&OKKK4YZJeRUMOIe77<:4GRRA
[YK&ykkk4t{skxyieozj4GRRA
{ok&rijevgiqgmk4GRRA

ktzyz&Luxskx&yo
Vuxz&.
&&&&&&&&YKW[KTIK&@&yt&YZJeRUMOIe\KIZUX&.7&zu&7</A&33&Хфчслкфижшлсђуфчшђ
&&&&&&&&J&@&yt&YZJeRUMOIe\KIZUX&.7&zu&?/A&33&Иёыфкё&шцоййлцфи
&&&&&&&&LXKW&@&yt&YZJeRUMOIe\KIZUX&.7;&ju}tzu&6/A&33&Эжчшфшж&76d.38/&Йь
&&&&&&&&SGT[GReSUJK&@&yt&YZJeRUMOIA&33&Цщэуфп&цлмот&3&72&жишф&3&6
&&&&&&&&VG[YK&@&yt&YZJeRUMOIA&33&Хжщнж&3&74
&&&&&&&&IRQ&@&yt&YZJeRUMOIA&33&Шжршфиёп&чойужс&ч&клсошлсѕ
&&&&&&&&
&&&&&&&&GXXG_eYZXOTM7&@&u{z&gxxgeule7<ehzkoezvkA&33&Хлцижѕ&чшцфрж
&&&&&&&&GXXG_eYZXOTM8&@&u{z&gxxgeule7<ehzkoezvk&33&Ишфцжѕ&чшцфрж
&&&&&/A
ktj&LuxskxA

gxinyzkiz{xk&Hkng|yuxgr&ul&Luxskx&yo
&&&&oymtgr&ZKSVeYZXOTM7@&gxxgeule7<ehzkoezvk@C&
&&&&.(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(/A
&&&&&
&&&&oymtgr&ZKSVeYZXOTM8@&gxxgeule7<ehzkoezvk&@C
&&&&.(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(2
&&&&&(66766666(/A
&&&&&
&&&&&l{tizyut&ingxezuehzk
&&&&&33&Ъщурьоѕ&хцлфзцжнщлш&иыфкуфп&чотифс&и&рфк&ѓшфйф&чотифсж&и&чффшилшчшиоо&ч&шжзсоьлп&
&&&&&33&чотифсфи&IM&XUS&о&ифницжяжлш&хфсщэлууфл&нужэлуол4&Лчсо&шжрфйф&чотифсж&улш&и&шжзсоьл2
&&&&&33&шф&ифницжяжлш&нужэлуол&хцфзлсж
&&&&&.
&&&&&&&&in@&INGXGIZKX
&&&&&/
&&&&&xkz{xt&hzkezvk&yo
&&&&&hkmyt
&&&&&&&&&&&&yl&&in&C&-&-&znkt&xkz{xt&(66766666(A
&&&&&&&&&&&&kroyl&in&C&-2-&znkt&xkz{xt&(66767766(A
&&&&&&&&&&&&kroyl&in&C&-6-&znkt&xkz{xt&(66776666(A
&&&&&&&&&&&&kroyl&in&C&-7-&znkt&xkz{xt&(66776667(A
&&&&&&&&&&&&kroyl&in&C&-8-&znkt&xkz{xt&(66776676(A
&&&&&&&&&&&&kroyl&in&C&-9-&znkt&xkz{xt&(66776677(A
&&&&&&&&&&&&kroyl&in&C&-:-&znkt&xkz{xt&(66776766(A
&&&&&&&&&&&&kroyl&in&C&-;-&znkt&xkz{xt&(66776767(A
&&&&&&&&&&&&kroyl&in&C&-<-&znkt&xkz{xt&(66776776(A
&&&&&&&&&&&&kroyl&in&C&-=-&znkt&xkz{xt&(66776777(A
&&&&&&&&&&&&kroyl&in&C&->-&znkt&xkz{xt&(66777666(A
&&&&&&&&&&&&kroyl&in&C&-?-&znkt&xkz{xt&(66777667(A
&&&&&&&&&&&&kroyl&in&C&-G-&znkt&xkz{xt&(67666667(A
&&&&&&&&&&&&kroyl&in&C&-H-&znkt&xkz{xt&(67666676(A
&&&&&&&&&&&&kroyl&in&C&-I-&znkt&xkz{xt&(67666677(A
&&&&&&&&&&&&kroyl&in&C&-J-&znkt&xkz{xt&(67666766(A
&&&&&&&&&&&&kroyl&in&C&-K-&znkt&xkz{xt&(67666767(A
&&&&&&&&&&&&kroyl&in&C&-L-&znkt&xkz{xt&(67666776(A
&&&&&&&&&&&&kroyl&in&C&-M-&znkt&xkz{xt&(67666777(A
&&&&&&&&&&&&kroyl&in&C&-N-&znkt&xkz{xt&(67667666(A
&&&&&&&&&&&&kroyl&in&C&-O-&znkt&xkz{xt&(67667667(A
&&&&&&&&&&&&kroyl&in&C&-P-&znkt&xkz{xt&(67667676(A
&&&&&&&&&&&&kroyl&in&C&-Q-&znkt&xkz{xt&(67667677(A
&&&&&&&&&&&&kroyl&in&C&-R-&znkt&xkz{xt&(67667766(A
&&&&&&&&&&&&kroyl&in&C&-S-&znkt&xkz{xt&(67667767(A
&&&&&&&&&&&&kroyl&in&C&-T-&znkt&xkz{xt&(67667776(A
&&&&&&&&&&&&kroyl&in&C&-U-&znkt&xkz{xt&(67667777(A
&&&&&&&&&&&&kroyl&in&C&-V-&znkt&xkz{xt&(67676666(A
&&&&&&&&&&&&kroyl&in&C&-W-&znkt&xkz{xt&(67676667(A
&&&&&&&&&&&&kroyl&in&C&-X-&znkt&xkz{xt&(67676676(A
&&&&&&&&&&&&kroyl&in&C&-Y-&znkt&xkz{xt&(67676677(A
&&&&&&&&&&&&kroyl&in&C&-Z-&znkt&xkz{xt&(67676766(A
&&&&&&&&&&&&kroyl&in&C&-[-&znkt&xkz{xt&(67676767(A
&&&&&&&&&&&&kroyl&in&C&-\-&znkt&xkz{xt&(67676776(A
&&&&&&&&&&&&kroyl&in&C&-]-&znkt&xkz{xt&(67676777(A
&&&&&&&&&&&&kroyl&in&C&-^-&znkt&xkz{xt&(67677666(A
&&&&&&&&&&&&kroyl&in&C&-_-&znkt&xkz{xt&(67677667(A
&&&&&&&&&&&&kroyl&in&C&-`-&znkt&xkz{xt&(67677676(A
&&&&&&&&&&&&krok&xkz{xt&(66766666(A
&&&&&&&&&&&&ktj&ylA
&&&&&ktj&ingxezuehzkA
&&&&
hkmyt
&&&&vxuikoo&.IRQ/&hkmyt
&&&&&&&&33&Нжхочђ&и&зщълцё&чшцфр&хф&ъцфушщ&отхщсђчж
&&&&&&&&yl&xyoytmekjmk.IRQ/&znkt
&&&&&&&&
&&&&&&&&&&&&33&Нжхочђ&зщълцж&хлцифп&чшцфро
&&&&&&&&&&&&R7@&lux&itz&yt&7&zu&7<&ruuv
&&&&&&&&&&&&&&&&yl&YKW[KTIK.itz/&C&-7-&znkt
&&&&&&&&&&&&&&&&&&&&ZKSVeYZXOTM7.itz/&BC&ingxezuehzk.-7-/A
&&&&&&&&&&&&&&&&krok
&&&&&&&&&&&&&&&&&&&&ZKSVeYZXOTM7.itz/&BC&ingxezuehzk.-6-/A
&&&&&&&&&&&&&&&&ktj&ylA
&&&&&&&&&&&&ktj&ruuv&R7A
&&&&&&&&&&&&
&&&&&&&&&&&&33&Нжхочђ&зщълцж&ишфцфп&чшфро&.чотифсё&7&3&?/
&&&&&&&&&&&&R8@&lux&itz&yt&7&zu&?&ruuv
&&&&&&&&&&&&&&&&yl&J.itz/&C&-7-&znkt
&&&&&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.itz/&BC&ingxezuehzk.-7-/A
&&&&&&&&&&&&&&&&kroyl&J.itz/&C&-6-&znkt
&&&&&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.itz/&BC&ingxezuehzk.-6-/A
&&&&&&&&&&&&&&&&krok
&&&&&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.itz/&BC&ingxezuehzk.-&-/A
&&&&&&&&&&&&&&&&ktj&ylA
&&&&&&&&&&&&ktj&ruuv&R8A
&&&&&&&&&&&&
&&&&&&&&ktj&ylA&
&&&&ktj&vxuikooA
&&&&
&&&&33&Нжхочђ&76фйф&чотифсж&ишфцфп&чшцфро
&&&&ZKSVeYZXOTM8.76/&BC&&(66666667(&]NKT&IRQ&C&-7-&KRYK
&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&(66666666(A
&&&&
&&&&vxuikoo&.SGT[GReSUJK2&VG[YK2&LXKW/
&&&&&&&&|gxyghrk&ZKSVeLXKW&@&ytzkmkx&xgtmk&6&zu&98=<>A
&&&&&&&&|gxyghrk&YZXOTMeLXKW&@&YZXOTM&.7&zu&;/A
&&&&&&&&hkmyt
&&&&&&&&
&&&&&&&&yl&VG[YK&C&-7-&znkt
&&&&&&&&&&&&ZKSVeYZXOTM8.77/&BC&ingxezuehzk.-V-/A
&&&&&&&&&&&&ZKSVeYZXOTM8.78/&BC&ingxezuehzk.-G-/A
&&&&&&&&&&&&ZKSVeYZXOTM8.79/&BC&ingxezuehzk.-[-/A
&&&&&&&&&&&&ZKSVeYZXOTM8.7:/&BC&ingxezuehzk.-Y-/A
&&&&&&&&&&&&ZKSVeYZXOTM8.7;/&BC&ingxezuehzk.-K-/A
&&&&&&&&&&&&ZKSVeYZXOTM8.7</&BC&ingxezuehzk.-&-/A
&&&&&&&&krok
&&&&&&&&&&&&yl&SGT[GReSUJK&C&-7-&znkt
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.77/&BC&ingxezuehzk.-S-/A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.78/&BC&ingxezuehzk.-G-/A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.79/&BC&ingxezuehzk.-T-/A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.7:/&BC&ingxezuehzk.-[-/A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.7;/&BC&ingxezuehzk.-G-/A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.7</&BC&ingxezuehzk.-R-/A
&&&&&&&&&&&&krok
&&&&&&&&&&&&&&&&ZKSVeLXKW&@C&ZUeOTZKMKX.[TYOMTKJ.LXKW//A
&&&&&&&&&&&&&&&&YZXOTMeLXKW&@C&ytzkmkx-ysgmk.ZKSVeLXKW/A

&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.77/&BC&ingxezuehzk.YZXOTMeLXKW.8//A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.78/&BC&ingxezuehzk.YZXOTMeLXKW.9//A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.79/&BC&ingxezuehzk.-2-/A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.7:/&BC&ingxezuehzk.YZXOTMeLXKW.://A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.7;/&BC&ingxezuehzk.YZXOTMeLXKW.;//A
&&&&&&&&&&&&&&&&ZKSVeYZXOTM8.7</&BC&(66666676(A&33&-N`-
&&&&&&&&&&&&ktj&ylA
&&&&&&&&ktj&ylA
&&&&ktj&vxuikooA
&&&&
&&&&GXXG_eYZXOTM7&BC&ZKSVeYZXOTM7A
&&&&GXXG_eYZXOTM8&BC&ZKSVeYZXOTM8A
&&&&
ktj&Hkng|yuxgrA
